module register65(out, in, clk, en, clr);
	input clk, en, clr;
	input signed [64:0] in;
	output signed [64:0] out;

	dffe_ref dfffe_0(out[0], in[0], clk, en, clr);
	dffe_ref dfffe_1(out[1], in[1], clk, en, clr);
	dffe_ref dfffe_2(out[2], in[2], clk, en, clr);
	dffe_ref dfffe_3(out[3], in[3], clk, en, clr);
	dffe_ref dfffe_4(out[4], in[4], clk, en, clr);
	dffe_ref dfffe_5(out[5], in[5], clk, en, clr);
	dffe_ref dfffe_6(out[6], in[6], clk, en, clr);
	dffe_ref dfffe_7(out[7], in[7], clk, en, clr);
	dffe_ref dfffe_8(out[8], in[8], clk, en, clr);
	dffe_ref dfffe_9(out[9], in[9], clk, en, clr);
	dffe_ref dfffe_10(out[10], in[10], clk, en, clr);
	dffe_ref dfffe_11(out[11], in[11], clk, en, clr);
	dffe_ref dfffe_12(out[12], in[12], clk, en, clr);
	dffe_ref dfffe_13(out[13], in[13], clk, en, clr);
	dffe_ref dfffe_14(out[14], in[14], clk, en, clr);
	dffe_ref dfffe_15(out[15], in[15], clk, en, clr);
	dffe_ref dfffe_16(out[16], in[16], clk, en, clr);
	dffe_ref dfffe_17(out[17], in[17], clk, en, clr);
	dffe_ref dfffe_18(out[18], in[18], clk, en, clr);
	dffe_ref dfffe_19(out[19], in[19], clk, en, clr);
	dffe_ref dfffe_20(out[20], in[20], clk, en, clr);
	dffe_ref dfffe_21(out[21], in[21], clk, en, clr);
	dffe_ref dfffe_22(out[22], in[22], clk, en, clr);
	dffe_ref dfffe_23(out[23], in[23], clk, en, clr);
	dffe_ref dfffe_24(out[24], in[24], clk, en, clr);
	dffe_ref dfffe_25(out[25], in[25], clk, en, clr);
	dffe_ref dfffe_26(out[26], in[26], clk, en, clr);
	dffe_ref dfffe_27(out[27], in[27], clk, en, clr);
	dffe_ref dfffe_28(out[28], in[28], clk, en, clr);
	dffe_ref dfffe_29(out[29], in[29], clk, en, clr);
	dffe_ref dfffe_30(out[30], in[30], clk, en, clr);
	dffe_ref dfffe_31(out[31], in[31], clk, en, clr);
	dffe_ref dfffe_32(out[32], in[32], clk, en, clr);
	dffe_ref dfffe_33(out[33], in[33], clk, en, clr);
	dffe_ref dfffe_34(out[34], in[34], clk, en, clr);
	dffe_ref dfffe_35(out[35], in[35], clk, en, clr);
	dffe_ref dfffe_36(out[36], in[36], clk, en, clr);
	dffe_ref dfffe_37(out[37], in[37], clk, en, clr);
	dffe_ref dfffe_38(out[38], in[38], clk, en, clr);
	dffe_ref dfffe_39(out[39], in[39], clk, en, clr);
	dffe_ref dfffe_40(out[40], in[40], clk, en, clr);
	dffe_ref dfffe_41(out[41], in[41], clk, en, clr);
	dffe_ref dfffe_42(out[42], in[42], clk, en, clr);
	dffe_ref dfffe_43(out[43], in[43], clk, en, clr);
	dffe_ref dfffe_44(out[44], in[44], clk, en, clr);
	dffe_ref dfffe_45(out[45], in[45], clk, en, clr);
	dffe_ref dfffe_46(out[46], in[46], clk, en, clr);
	dffe_ref dfffe_47(out[47], in[47], clk, en, clr);
	dffe_ref dfffe_48(out[48], in[48], clk, en, clr);
	dffe_ref dfffe_49(out[49], in[49], clk, en, clr);
	dffe_ref dfffe_50(out[50], in[50], clk, en, clr);
	dffe_ref dfffe_51(out[51], in[51], clk, en, clr);
	dffe_ref dfffe_52(out[52], in[52], clk, en, clr);
	dffe_ref dfffe_53(out[53], in[53], clk, en, clr);
	dffe_ref dfffe_54(out[54], in[54], clk, en, clr);
	dffe_ref dfffe_55(out[55], in[55], clk, en, clr);
	dffe_ref dfffe_56(out[56], in[56], clk, en, clr);
	dffe_ref dfffe_57(out[57], in[57], clk, en, clr);
	dffe_ref dfffe_58(out[58], in[58], clk, en, clr);
	dffe_ref dfffe_59(out[59], in[59], clk, en, clr);
	dffe_ref dfffe_60(out[60], in[60], clk, en, clr);
	dffe_ref dfffe_61(out[61], in[61], clk, en, clr);
	dffe_ref dfffe_62(out[62], in[62], clk, en, clr);
	dffe_ref dfffe_63(out[63], in[63], clk, en, clr);
	dffe_ref dfffe_64(out[64], in[64], clk, en, clr);
endmodule
