module not32(data_result, data_operandA);
        
    input [31:0] data_operandA;

    output [31:0] data_result;

    not bit0 (data_result[0], data_operandA[0]);
    not bit1 (data_result[1], data_operandA[1]);
    not bit2 (data_result[2], data_operandA[2]);
    not bit3 (data_result[3], data_operandA[3]);
    not bit4 (data_result[4], data_operandA[4]);
    not bit5 (data_result[5], data_operandA[5]);
    not bit6 (data_result[6], data_operandA[6]);
    not bit7 (data_result[7], data_operandA[7]);
    not bit8 (data_result[8], data_operandA[8]);
    not bit9 (data_result[9], data_operandA[9]);
    not bit10 (data_result[10], data_operandA[10]);
    not bit11 (data_result[11], data_operandA[11]);
    not bit12 (data_result[12], data_operandA[12]);
    not bit13 (data_result[13], data_operandA[13]);
    not bit14 (data_result[14], data_operandA[14]);
    not bit15 (data_result[15], data_operandA[15]);
    not bit16 (data_result[16], data_operandA[16]);
    not bit17 (data_result[17], data_operandA[17]);
    not bit18 (data_result[18], data_operandA[18]);
    not bit19 (data_result[19], data_operandA[19]);
    not bit20 (data_result[20], data_operandA[20]);
    not bit21 (data_result[21], data_operandA[21]);
    not bit22 (data_result[22], data_operandA[22]);
    not bit23 (data_result[23], data_operandA[23]);
    not bit24 (data_result[24], data_operandA[24]);
    not bit25 (data_result[25], data_operandA[25]);
    not bit26 (data_result[26], data_operandA[26]);
    not bit27 (data_result[27], data_operandA[27]);
    not bit28 (data_result[28], data_operandA[28]);
    not bit29 (data_result[29], data_operandA[29]);
    not bit30 (data_result[30], data_operandA[30]);
    not bit31 (data_result[31], data_operandA[31]);

endmodule